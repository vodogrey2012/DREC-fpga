
module unnamed (
	noe_in);	

	input		noe_in;
endmodule
