// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// Created on Fri Nov  5 18:47:12 2021

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    reset,clock,btn1,btn2,btn4,
    led1,led2);

    input reset;
    input clock;
    input btn1;
    input btn2;
    input btn4;
    tri0 reset;
    tri0 btn1;
    tri0 btn2;
    tri0 btn4;
    output led1;
    output led2;
    reg led1;
    reg led2;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or btn1 or btn2 or btn4)
    begin
        if (reset) begin
            reg_fstate <= state1;
            led1 <= 1'b0;
            led2 <= 1'b0;
        end
        else begin
            led1 <= 1'b0;
            led2 <= 1'b0;
            case (fstate)
                state1: begin
                    if (~(btn1))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    led1 <= 1'b1;

                    led2 <= 1'b1;
                end
                state2: begin
                    if ((~(btn2) & btn4))
                        reg_fstate <= state3;
                    else if ((~(btn4) & btn2))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    led1 <= 1'b0;

                    led2 <= 1'b1;
                end
                state3: begin
                    if ((~(btn1) & btn4))
                        reg_fstate <= state4;
                    else if ((~(btn4) & btn1))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    led1 <= 1'b1;

                    led2 <= 1'b0;
                end
                state4: begin
                    if ((~(btn2) | ~(btn4)))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    led1 <= 1'b0;

                    led2 <= 1'b0;
                end
                default: begin
                    led1 <= 1'bx;
                    led2 <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM1
